LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
USE IEEE.numeric_std.ALL;

ENTITY FIR32_DecimateBy2_abstracted IS
    PORT( 
        clk_Fs_x8       :   IN    std_logic;  -- system clock rate: Fs times 8 (due to folding)
        clk_Fs          :   IN    std_logic;  -- input  clock rate: Fs
        clk_Fs_d2       :   IN    std_logic;  -- output clock rate: Fs divided by 2
        reset           :   IN    std_logic;
        data_in         :   IN    std_logic_vector(31 DOWNTO 0); -- sfix32_En28  -- data in  at Fs   rate
        data_out        :   OUT   std_logic_vector(31 DOWNTO 0)  -- sfix32_En28  -- data out at Fs/2 rate
    );
END FIR32_DecimateBy2_abstracted;


ARCHITECTURE rtl OF FIR32_DecimateBy2_abstracted IS

    component FIR32_DecimateBy2 IS
       PORT( clk                             :   IN    std_logic; 
             clk_enable                      :   IN    std_logic; 
             reset                           :   IN    std_logic; 
             filter_in                       :   IN    std_logic_vector(31 DOWNTO 0); -- sfix32_En28
             filter_out                      :   OUT   std_logic_vector(68 DOWNTO 0); -- sfix69_En60
             ce_out                          :   OUT   std_logic  
             );
    
    END component;
    --### Clock rate is 8 times the input and 16 times the output sample rate for this architecture.
    --### Successful completion of VHDL code generation process for filter: FIR32_DecimateBy2
    --### HDL latency is 2 samples
    -- Code auto generated by Matlab:  filter_length = 64; 
    --                            down_converter = dsp.FIRDecimator(2,fir1(filter_length,0.48));
    --                            fdhdltool(down_converter,numerictype(1,32,28))
    
 	-- decimator signals
	signal  decimator_data_in     : std_logic_vector(31 DOWNTO 0); -- sfix32_En28
	signal  decimator_data_out    : std_logic_vector(68 DOWNTO 0); -- sfix69_En60  
	signal  data_out_int          : std_logic_vector(68 DOWNTO 0); -- sfix69_En60   
	--signal  decimator_ce_out      : std_logic;   
	 
BEGIN

    -------------------------------------------------------------------
    -- Capture data in on Fs clock
    -------------------------------------------------------------------
    process(clk_Fs)
    begin
        if rising_edge(clk_Fs) then
            decimator_data_in <= data_in;
        end if;
    end process;
    
    -------------------------------------------------------------------
    -- Send through decimator
    -------------------------------------------------------------------
	decimator : FIR32_DecimateBy2 port map (
		clk         =>  clk_Fs_x8,                       
		clk_enable  =>  '1',
		reset       =>  reset,
		filter_in   =>  decimator_data_in,      
		filter_out  =>  decimator_data_out,
		ce_out      =>  open
	);
     
     
    -------------------------------------------------------------------
    -- output data on Fs/2 clock
    -------------------------------------------------------------------
    process(clk_Fs_d2)
    begin
        if rising_edge(clk_Fs_d2) then   
            data_out <= decimator_data_out(63 downto 32);  -- convert back to -- sfix32_En28
        end if;
    end process;
     

END rtl;