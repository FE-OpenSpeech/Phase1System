LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
USE IEEE.numeric_std.ALL;

ENTITY FIR32_InterpolateBy2_abstracted IS
    PORT( 
        clk_Fs_x16      :   IN    std_logic;  -- system clock rate: Fs times 32 (due to folding)
        clk_Fs          :   IN    std_logic;  -- input  clock rate: Fs
        clk_Fs_x2       :   IN    std_logic;  -- output clock rate: Fs times 2
        reset           :   IN    std_logic;
        data_in         :   IN    std_logic_vector(31 DOWNTO 0); -- sfix32_En28  -- data in  at Fs   rate
        data_out        :   OUT   std_logic_vector(31 DOWNTO 0)  -- sfix32_En28  -- data out at Fs*2 rate
    );
END FIR32_InterpolateBy2_abstracted;


ARCHITECTURE rtl OF FIR32_InterpolateBy2_abstracted IS

    component FIR32_InterpolateBy2 IS
       PORT( clk                             :   IN    std_logic; 
             clk_enable                      :   IN    std_logic; 
             reset                           :   IN    std_logic; 
             filter_in                       :   IN    std_logic_vector(31 DOWNTO 0); -- sfix32_En28
             filter_out                      :   OUT   std_logic_vector(68 DOWNTO 0); -- sfix70_En60
             ce_out                          :   OUT   std_logic  
             );
    
    END component;
    --### Clock rate is 16 times the input and 8 times the output sample rate for this architecture.
    --### Successful completion of VHDL code generation process for filter: FIR32_InterpolateBy2
    --### HDL latency is 1 samples
    -- Code auto generated by Matlab:  filter_length = 32; 
    --                            up_converter = dsp.FIRInterpolator(2,fir1(filter_length,0.48));
    --                            fdhdltool(up_converter,numerictype(1,32,28))
    
 	-- interpolator signals
	signal  interpolator_data_in  : std_logic_vector(31 DOWNTO 0); -- sfix32_En28
	signal  interpolator_data_out : std_logic_vector(68 DOWNTO 0); -- sfix70_En60  
	signal  data_out_int          : std_logic_vector(68 DOWNTO 0); -- sfix70_En60   
	--signal  interpolator_ce_out   : std_logic;   
	 
BEGIN

    -------------------------------------------------------------------
    -- Capture data in on Fs clock
    -------------------------------------------------------------------
    process(clk_Fs)
    begin
        if rising_edge(clk_Fs) then
            interpolator_data_in <= data_in;
        end if;
    end process;
    
    -------------------------------------------------------------------
    -- Send through interpolator
    -------------------------------------------------------------------
	interpolator : FIR32_InterpolateBy2 port map (
		clk         =>  clk_Fs_x16,                       
		clk_enable  =>  '1',
		reset       =>  reset,
		filter_in   =>  interpolator_data_in,      
		filter_out  =>  interpolator_data_out,
		ce_out      =>  open
	);
          
    -------------------------------------------------------------------
    -- output data on Fs*2 clock
    -------------------------------------------------------------------
    process(clk_Fs_x2)
    begin
        if rising_edge(clk_Fs_x2) then   
            data_out <= interpolator_data_out(62 downto 31);  -- convert back to -- sfix32_En28
        end if;
    end process;
     

END rtl;